`include "axi_interface.sv"
`include "axi_transaction.sv"
`include "axi_sequencer.sv"
`include "axi_driver.sv"
`include "axi_monitor.sv"
`include "axi_agent.sv"
`include "axi_scoreboard.sv"
`include "axi_subscriber.sv"
`include "axi_environment.sv"
`include "axi_sequence.sv"
`include "axi_test.sv"