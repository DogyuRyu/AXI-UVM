module axi_interface_adapter #(
  parameter AXI_DW = 64,
  parameter AXI_AW = 32,
  parameter AXI_IW = 8,
  parameter AXI_SW = AXI_DW/8
)(
  // AXI4 인터페이스 (BFM 쪽)
  AXI4 #(.N(AXI_SW), .I(AXI_IW)) bfm_intf,
  
  // AXI3 신호 (DUT 쪽)
  // global signals
  output                    axi_clk_i,
  output                    axi_rstn_i,
  
  // axi write address channel
  output     [ AXI_IW-1: 0] axi_awid_i,
  output     [ AXI_AW-1: 0] axi_awaddr_i,
  output     [      4-1: 0] axi_awlen_i,  // AXI3는 4비트 AWLEN
  output     [      3-1: 0] axi_awsize_i,
  output     [      2-1: 0] axi_awburst_i,
  output     [      2-1: 0] axi_awlock_i,
  output     [      4-1: 0] axi_awcache_i,
  output     [      3-1: 0] axi_awprot_i,
  output                    axi_awvalid_i,
  input                     axi_awready_o,
  
  // axi write data channel
  output     [ AXI_IW-1: 0] axi_wid_i,    // AXI3에는 WID 존재
  output     [ AXI_DW-1: 0] axi_wdata_i,
  output     [ AXI_SW-1: 0] axi_wstrb_i,
  output                    axi_wlast_i,
  output                    axi_wvalid_i,
  input                     axi_wready_o,
  
  // axi write response channel
  input      [ AXI_IW-1: 0] axi_bid_o,
  input      [      2-1: 0] axi_bresp_o,
  input                     axi_bvalid_o,
  output                    axi_bready_i,
  
  // axi read address channel
  output     [ AXI_IW-1: 0] axi_arid_i,
  output     [ AXI_AW-1: 0] axi_araddr_i,
  output     [      4-1: 0] axi_arlen_i,  // AXI3는 4비트 ARLEN
  output     [      3-1: 0] axi_arsize_i,
  output     [      2-1: 0] axi_arburst_i,
  output     [      2-1: 0] axi_arlock_i,
  output     [      4-1: 0] axi_arcache_i,
  output     [      3-1: 0] axi_arprot_i,
  output                    axi_arvalid_i,
  input                     axi_arready_o,
  
  // axi read data channel
  input      [ AXI_IW-1: 0] axi_rid_o,
  input      [ AXI_DW-1: 0] axi_rdata_o,
  input      [      2-1: 0] axi_rresp_o,
  input                     axi_rlast_o,
  input                     axi_rvalid_o,
  output                    axi_rready_i,
  
  // 시스템 버스 신호 (DUT 특화)
  input      [ AXI_AW-1: 0] sys_addr_o,
  input      [ AXI_DW-1: 0] sys_wdata_o,
  input      [ AXI_SW-1: 0] sys_sel_o,
  input                     sys_wen_o,
  input                     sys_ren_o,
  output     [ AXI_DW-1: 0] sys_rdata_i,
  output                    sys_err_i,
  output                    sys_ack_i
);

  // 클럭 및 리셋 연결
  assign axi_clk_i = bfm_intf.ACLK;
  assign axi_rstn_i = bfm_intf.ARESETn;
  
  // Write Address 채널 연결
  assign axi_awid_i = bfm_intf.AWID;
  assign axi_awaddr_i = bfm_intf.AWADDR;
  assign axi_awlen_i = bfm_intf.AWLEN[3:0]; // AXI4 -> AXI3 변환
  assign axi_awsize_i = bfm_intf.AWSIZE;
  assign axi_awburst_i = bfm_intf.AWBURST;
  assign axi_awlock_i = {1'b0, bfm_intf.AWLOCK}; // AXI4는 1비트, AXI3는 2비트
  assign axi_awcache_i = bfm_intf.AWCACHE;
  assign axi_awprot_i = bfm_intf.AWPROT;
  assign axi_awvalid_i = bfm_intf.AWVALID;
  assign bfm_intf.AWREADY = axi_awready_o;
  
  // Write Data 채널 연결
  assign axi_wid_i = bfm_intf.AWID; // AXI4에는 WID가 없으므로 AWID 사용
  assign axi_wdata_i = bfm_intf.WDATA;
  assign axi_wstrb_i = bfm_intf.WSTRB;
  assign axi_wlast_i = bfm_intf.WLAST;
  assign axi_wvalid_i = bfm_intf.WVALID;
  assign bfm_intf.WREADY = axi_wready_o;
  
  // Write Response 채널 연결
  assign bfm_intf.BID = axi_bid_o;
  assign bfm_intf.BRESP = axi_bresp_o;
  assign bfm_intf.BVALID = axi_bvalid_o;
  assign axi_bready_i = bfm_intf.BREADY;
  
  // Read Address 채널 연결
  assign axi_arid_i = bfm_intf.ARID;
  assign axi_araddr_i = bfm_intf.ARADDR;
  assign axi_arlen_i = bfm_intf.ARLEN[3:0]; // AXI4 -> AXI3 변환
  assign axi_arsize_i = bfm_intf.ARSIZE;
  assign axi_arburst_i = bfm_intf.ARBURST;
  assign axi_arlock_i = {1'b0, bfm_intf.ARLOCK}; // AXI4는 1비트, AXI3는 2비트
  assign axi_arcache_i = bfm_intf.ARCACHE;
  assign axi_arprot_i = bfm_intf.ARPROT;
  assign axi_arvalid_i = bfm_intf.ARVALID;
  assign bfm_intf.ARREADY = axi_arready_o;
  
  // Read Data 채널 연결
  assign bfm_intf.RID = axi_rid_o;
  assign bfm_intf.RDATA = axi_rdata_o;
  assign bfm_intf.RRESP = axi_rresp_o;
  assign bfm_intf.RLAST = axi_rlast_o;
  assign bfm_intf.RVALID = axi_rvalid_o;
  assign axi_rready_i = bfm_intf.RREADY;
  
  // 시스템 버스 신호 (필요에 따라 연결)
  assign sys_rdata_i = 64'h0; // 기본값, 필요에 따라 변경
  assign sys_err_i = 1'b0;     // 기본값, 필요에 따라 변경
  assign sys_ack_i = 1'b1;     // 기본값, 필요에 따라 변경
  
endmodule