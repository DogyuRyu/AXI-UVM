`include "interface.sv"
`include "transaction.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "subscriber.sv"
`include "environment.sv"
`include "sequence.sv"
`include "test.sv"